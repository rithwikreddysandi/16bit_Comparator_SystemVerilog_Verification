// Transaction Class

class comp_tx;
  rand bit [15:0] a,b; // randomizing the a,b to compare these 16-bit inputs
  bit [0:0]  less, equal, greater;
endclass